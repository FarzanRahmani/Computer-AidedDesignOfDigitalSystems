library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.Numeric_STD.ALL;

package types is 
	
	type array_of_8bit is array(0 to 9) of std_logic_vector(0 to 7);

	
end types;